module SubByte (input [7:0] State,output reg [7:0] Statep);

always @(State)


case(State)

8'h00: Statep=8'h63;
8'h01: Statep=8'h7c;
8'h02: Statep=8'h77;
8'h03: Statep=8'h7b;
8'h04: Statep=8'hf2;
8'h05: Statep=8'h6b;
8'h06: Statep=8'h6f;
8'h07: Statep=8'hc5;
8'h08: Statep=8'h30;
8'h09: Statep=8'h01;
8'h0a: Statep=8'h67;
8'h0b: Statep=8'h2b;
8'h0c: Statep=8'hfe;
8'h0d: Statep=8'hd7;
8'h0e: Statep=8'hab;
8'h0f: Statep=8'h76;
8'h10: Statep=8'hca;
8'h11: Statep=8'h82;
8'h12: Statep=8'hc9;
8'h13: Statep=8'h7d;
8'h14: Statep=8'hfa;
8'h15: Statep=8'h59;
8'h16: Statep=8'h47;
8'h17: Statep=8'hf0;
8'h18: Statep=8'had;
8'h19: Statep=8'hd4;
8'h1a: Statep=8'ha2;
8'h1b: Statep=8'haf;
8'h1c: Statep=8'h9c;
8'h1d: Statep=8'ha4;
8'h1e: Statep=8'h72;
8'h1f: Statep=8'hc0;
8'h20: Statep=8'hb7;
8'h21: Statep=8'hfd;
8'h22: Statep=8'h93;
8'h23: Statep=8'h26;
8'h24: Statep=8'h36;
8'h25: Statep=8'h3f;
8'h26: Statep=8'hf7;
8'h27: Statep=8'hcc;
8'h28: Statep=8'h34;
8'h29: Statep=8'ha5;
8'h2a: Statep=8'he5;
8'h2b: Statep=8'hf1;
8'h2c: Statep=8'h71;
8'h2d: Statep=8'hd8;
8'h2e: Statep=8'h31;
8'h2f: Statep=8'h15;
8'h30: Statep=8'h04;
8'h31: Statep=8'hc7;
8'h32: Statep=8'h23;
8'h33: Statep=8'hc3;
8'h34: Statep=8'h18;
8'h35: Statep=8'h96;
8'h36: Statep=8'h05;
8'h37: Statep=8'h9a;
8'h38: Statep=8'h07;
8'h39: Statep=8'h12;
8'h3a: Statep=8'h80;
8'h3b: Statep=8'he2;
8'h3c: Statep=8'heb;
8'h3d: Statep=8'h27;
8'h3e: Statep=8'hb2;
8'h3f: Statep=8'h75;
8'h40: Statep=8'h09;
8'h41: Statep=8'h83;
8'h42: Statep=8'h2c;
8'h43: Statep=8'h1a;
8'h44: Statep=8'h1b;
8'h45: Statep=8'h6e;
8'h46: Statep=8'h5a;
8'h47: Statep=8'ha0;
8'h48: Statep=8'h52;
8'h49: Statep=8'h3b;
8'h4a: Statep=8'hd6;
8'h4b: Statep=8'hb3;
8'h4c: Statep=8'h29;
8'h4d: Statep=8'he3;
8'h4e: Statep=8'h2f;
8'h4f: Statep=8'h84;
8'h50: Statep=8'h53;
8'h51: Statep=8'hd1;
8'h52: Statep=8'h00;
8'h53: Statep=8'hed;
8'h54: Statep=8'h20;
8'h55: Statep=8'hfc;
8'h56: Statep=8'hb1;
8'h57: Statep=8'h5b;
8'h58: Statep=8'h6a;
8'h59: Statep=8'hcb;
8'h5a: Statep=8'hbe;
8'h5b: Statep=8'h39;
8'h5c: Statep=8'h4a;
8'h5d: Statep=8'h4c;
8'h5e: Statep=8'h58;
8'h5f: Statep=8'hcf;
8'h60: Statep=8'hd0;
8'h61: Statep=8'hef;
8'h62: Statep=8'haa;
8'h63: Statep=8'hfb;
8'h64: Statep=8'h43;
8'h65: Statep=8'h4d;
8'h66: Statep=8'h33;
8'h67: Statep=8'h85;
8'h68: Statep=8'h45;
8'h69: Statep=8'hf9;
8'h6a: Statep=8'h02;
8'h6b: Statep=8'h7f;
8'h6c: Statep=8'h50;
8'h6d: Statep=8'h3c;
8'h6e: Statep=8'h9f;
8'h6f: Statep=8'ha8;
8'h70: Statep=8'h51;
8'h71: Statep=8'ha3;
8'h72: Statep=8'h40;
8'h73: Statep=8'h8f;
8'h74: Statep=8'h92;
8'h75: Statep=8'h9d;
8'h76: Statep=8'h38;
8'h77: Statep=8'hf5;
8'h78: Statep=8'hbc;
8'h79: Statep=8'hb6;
8'h7a: Statep=8'hda;
8'h7b: Statep=8'h21;
8'h7c: Statep=8'h10;
8'h7d: Statep=8'hff;
8'h7e: Statep=8'hf3;
8'h7f: Statep=8'hd2;
8'h80: Statep=8'hcd;
8'h81: Statep=8'h0c;
8'h82: Statep=8'h13;
8'h83: Statep=8'hec;
8'h84: Statep=8'h5f;
8'h85: Statep=8'h97;
8'h86: Statep=8'h44;
8'h87: Statep=8'h17;
8'h88: Statep=8'hc4;
8'h89: Statep=8'ha7;
8'h8a: Statep=8'h7e;
8'h8b: Statep=8'h3d;
8'h8c: Statep=8'h64;
8'h8d: Statep=8'h5d;
8'h8e: Statep=8'h19;
8'h8f: Statep=8'h73;
8'h90: Statep=8'h60;
8'h91: Statep=8'h81;
8'h92: Statep=8'h4f;
8'h93: Statep=8'hdc;
8'h94: Statep=8'h22;
8'h95: Statep=8'h2a;
8'h96: Statep=8'h90;
8'h97: Statep=8'h88;
8'h98: Statep=8'h46;
8'h99: Statep=8'hee;
8'h9a: Statep=8'hb8;
8'h9b: Statep=8'h14;
8'h9c: Statep=8'hde;
8'h9d: Statep=8'h5e;
8'h9e: Statep=8'h0b;
8'h9f: Statep=8'hdb;
8'ha0: Statep=8'he0;
8'ha1: Statep=8'h32;
8'ha2: Statep=8'h3a;
8'ha3: Statep=8'h0a;
8'ha4: Statep=8'h49;
8'ha5: Statep=8'h06;
8'ha6: Statep=8'h24;
8'ha7: Statep=8'h5c;
8'ha8: Statep=8'hc2;
8'ha9: Statep=8'hd3;
8'haa: Statep=8'hac;
8'hab: Statep=8'h62;
8'hac: Statep=8'h91;
8'had: Statep=8'h95;
8'hae: Statep=8'he4;
8'haf: Statep=8'h79;
8'hb0: Statep=8'he7;
8'hb1: Statep=8'hc8;
8'hb2: Statep=8'h37;
8'hb3: Statep=8'h6d;
8'hb4: Statep=8'h8d;
8'hb5: Statep=8'hd5;
8'hb6: Statep=8'h4e;
8'hb7: Statep=8'ha9;
8'hb8: Statep=8'h6c;
8'hb9: Statep=8'h56;
8'hba: Statep=8'hf4;
8'hbb: Statep=8'hea;
8'hbc: Statep=8'h65;
8'hbd: Statep=8'h7a;
8'hbe: Statep=8'hae;
8'hbf: Statep=8'h08;
8'hc0: Statep=8'hba;
8'hc1: Statep=8'h78;
8'hc2: Statep=8'h25;
8'hc3: Statep=8'h2e;
8'hc4: Statep=8'h1c;
8'hc5: Statep=8'ha6;
8'hc6: Statep=8'hb4;
8'hc7: Statep=8'hc6;
8'hc8: Statep=8'he8;
8'hc9: Statep=8'hdd;
8'hca: Statep=8'h74;
8'hcb: Statep=8'h1f;
8'hcc: Statep=8'h4b;
8'hcd: Statep=8'hbd;
8'hce: Statep=8'h8b;
8'hcf: Statep=8'h8a;
8'hd0: Statep=8'h70;
8'hd1: Statep=8'h3e;
8'hd2: Statep=8'hb5;
8'hd3: Statep=8'h66;
8'hd4: Statep=8'h48;
8'hd5: Statep=8'h03;
8'hd6: Statep=8'hf6;
8'hd7: Statep=8'h0e;
8'hd8: Statep=8'h61;
8'hd9: Statep=8'h35;
8'hda: Statep=8'h57;
8'hdb: Statep=8'hb9;
8'hdc: Statep=8'h86;
8'hdd: Statep=8'hc1;
8'hde: Statep=8'h1d;
8'hdf: Statep=8'h9e;
8'he0: Statep=8'he1;
8'he1: Statep=8'hf8;
8'he2: Statep=8'h98;
8'he3: Statep=8'h11;
8'he4: Statep=8'h69;
8'he5: Statep=8'hd9;
8'he6: Statep=8'h8e;
8'he7: Statep=8'h94;
8'he8: Statep=8'h9b;
8'he9: Statep=8'h1e;
8'hea: Statep=8'h87;
8'heb: Statep=8'he9;
8'hec: Statep=8'hce;
8'hed: Statep=8'h55;
8'hee: Statep=8'h28;
8'hef: Statep=8'hdf;
8'hf0: Statep=8'h8c;
8'hf1: Statep=8'ha1;
8'hf2: Statep=8'h89;
8'hf3: Statep=8'h0d;
8'hf4: Statep=8'hbf;
8'hf5: Statep=8'he6;
8'hf6: Statep=8'h42;
8'hf7: Statep=8'h68;
8'hf8: Statep=8'h41;
8'hf9: Statep=8'h99;
8'hfa: Statep=8'h2d;
8'hfb: Statep=8'h0f;
8'hfc: Statep=8'hb0;
8'hfd: Statep=8'h54;
8'hfe: Statep=8'hbb;
8'hff: Statep=8'h16;

endcase

endmodule