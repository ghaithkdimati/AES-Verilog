module InvSubBytes(state,nextstate);
input [0:7] state;
output [0:7] nextstate;
reg [0:7] tempout;
assign nextstate=tempout;
always @*
begin 
case(state)
8'h00: tempout=8'h52;
8'h01: tempout=8'h09;
8'h02: tempout=8'h6a;
8'h03: tempout=8'hd5;
8'h04: tempout=8'h30;
8'h05: tempout=8'h36;
8'h06: tempout=8'ha5;
8'h07: tempout=8'h38;
8'h08: tempout=8'hbf;
8'h09: tempout=8'h40;
8'h0a: tempout=8'ha3;
8'h0b: tempout=8'h9e;
8'h0c: tempout=8'h81;
8'h0d: tempout=8'hf3;
8'h0e: tempout=8'hd7;
8'h0f: tempout=8'hfb;
8'h10: tempout=8'h7c;
8'h11: tempout=8'he3;
8'h12: tempout=8'h39;
8'h13: tempout=8'h82;
8'h14: tempout=8'h9b;
8'h15: tempout=8'h2f;
8'h16: tempout=8'hff;
8'h17: tempout=8'h87;
8'h18: tempout=8'h34;
8'h19: tempout=8'h8e;
8'h1a: tempout=8'h43;
8'h1b: tempout=8'h44;
8'h1c: tempout=8'hc4;
8'h1d: tempout=8'hde;
8'h1e: tempout=8'he9;
8'h1f: tempout=8'hcb;
8'h20: tempout=8'h54;
8'h21: tempout=8'h7b;
8'h22: tempout=8'h94;
8'h23: tempout=8'h32;
8'h24: tempout=8'ha6;
8'h25: tempout=8'hc2;
8'h26: tempout=8'h23;
8'h27: tempout=8'h3d;
8'h28: tempout=8'hee;
8'h29: tempout=8'h4c;
8'h2a: tempout=8'h95;
8'h2b: tempout=8'h0b;
8'h2c: tempout=8'h42;
8'h2d: tempout=8'hfa;
8'h2e: tempout=8'hc3;
8'h2f: tempout=8'h4e;
8'h30: tempout=8'h08;
8'h31: tempout=8'h2e;
8'h32: tempout=8'ha1;
8'h33: tempout=8'h66;
8'h34: tempout=8'h28;
8'h35: tempout=8'hd9;
8'h36: tempout=8'h24;
8'h37: tempout=8'hb2;
8'h38: tempout=8'h76;
8'h39: tempout=8'h5b;
8'h3a: tempout=8'ha2;
8'h3b: tempout=8'h49;
8'h3c: tempout=8'h6d;
8'h3d: tempout=8'h8b;
8'h3e: tempout=8'hd1;
8'h3f: tempout=8'h25;
8'h40: tempout=8'h72;
8'h41: tempout=8'hf8;
8'h42: tempout=8'hf6;
8'h43: tempout=8'h64;
8'h44: tempout=8'h86;
8'h45: tempout=8'h68;
8'h46: tempout=8'h98;
8'h47: tempout=8'h16;
8'h48: tempout=8'hd4;
8'h49: tempout=8'ha4;
8'h4a: tempout=8'h5c;
8'h4b: tempout=8'hcc;
8'h4c: tempout=8'h5d;
8'h4d: tempout=8'h65;
8'h4e: tempout=8'hb6;
8'h4f: tempout=8'h92;
8'h50: tempout=8'h6c;
8'h51: tempout=8'h70;
8'h52: tempout=8'h48;
8'h53: tempout=8'h50;
8'h54: tempout=8'hfd;
8'h55: tempout=8'hed;
8'h56: tempout=8'hb9;
8'h57: tempout=8'hda;
8'h58: tempout=8'h5e;
8'h59: tempout=8'h15;
8'h5a: tempout=8'h46;
8'h5b: tempout=8'h57;
8'h5c: tempout=8'ha7;
8'h5d: tempout=8'h8d;
8'h5e: tempout=8'h9d;
8'h5f: tempout=8'h84;
8'h60: tempout=8'h90;
8'h61: tempout=8'hd8;
8'h62: tempout=8'hab;
8'h63: tempout=8'h00;
8'h64: tempout=8'h8c;
8'h65: tempout=8'hbc;
8'h66: tempout=8'hd3;
8'h67: tempout=8'h0a;
8'h68: tempout=8'hf7;
8'h69: tempout=8'he4;
8'h6a: tempout=8'h58;
8'h6b: tempout=8'h05;
8'h6c: tempout=8'hb8;
8'h6d: tempout=8'hb3;
8'h6e: tempout=8'h45;
8'h6f: tempout=8'h06;
8'h70: tempout=8'hd0;
8'h71: tempout=8'h2c;
8'h72: tempout=8'h1e;
8'h73: tempout=8'h8f;
8'h74: tempout=8'hca;
8'h75: tempout=8'h3f;
8'h76: tempout=8'h0f;
8'h77: tempout=8'h02;
8'h78: tempout=8'hc1;
8'h79: tempout=8'haf;
8'h7a: tempout=8'hbd;
8'h7b: tempout=8'h03;
8'h7c: tempout=8'h01;
8'h7d: tempout=8'h13;
8'h7e: tempout=8'h8a;
8'h7f: tempout=8'h6b;
8'h80: tempout=8'h3a;
8'h81: tempout=8'h91;
8'h82: tempout=8'h11;
8'h83: tempout=8'h41;
8'h84: tempout=8'h4f;
8'h85: tempout=8'h67;
8'h86: tempout=8'hdc;
8'h87: tempout=8'hea;
8'h88: tempout=8'h97;
8'h89: tempout=8'hf2;
8'h8a: tempout=8'hcf;
8'h8b: tempout=8'hce;
8'h8c: tempout=8'hf0;
8'h8d: tempout=8'hb4;
8'h8e: tempout=8'he6;
8'h8f: tempout=8'h73;
8'h90: tempout=8'h96;
8'h91: tempout=8'hac;
8'h92: tempout=8'h74;
8'h93: tempout=8'h22;
8'h94: tempout=8'he7;
8'h95: tempout=8'had;
8'h96: tempout=8'h35;
8'h97: tempout=8'h85;
8'h98: tempout=8'he2;
8'h99: tempout=8'hf9;
8'h9a: tempout=8'h37;
8'h9b: tempout=8'he8;
8'h9c: tempout=8'h1c;
8'h9d: tempout=8'h75;
8'h9e: tempout=8'hdf;
8'h9f: tempout=8'h6e;
8'ha0: tempout=8'h47;
8'ha1: tempout=8'hf1;
8'ha2: tempout=8'h1a;
8'ha3: tempout=8'h71;
8'ha4: tempout=8'h1d;
8'ha5: tempout=8'h29;
8'ha6: tempout=8'hc5;
8'ha7: tempout=8'h89;
8'ha8: tempout=8'h6f;
8'ha9: tempout=8'hb7;
8'haa: tempout=8'h62;
8'hab: tempout=8'h0e;
8'hac: tempout=8'haa; 
8'had: tempout=8'h18;
8'hae: tempout=8'hbe;
8'haf: tempout=8'h1b;
8'hb0: tempout=8'hfc;
8'hb1: tempout=8'h56;
8'hb2: tempout=8'h3e;
8'hb3: tempout=8'h4b;
8'hb4: tempout=8'hc6;
8'hb5: tempout=8'hd2;
8'hb6: tempout=8'h79;
8'hb7: tempout=8'h20;
8'hb8: tempout=8'h9a;
8'hb9: tempout=8'hdb;
8'hba: tempout=8'hc0;
8'hbb: tempout=8'hfe;
8'hbc: tempout=8'h78;
8'hbd: tempout=8'hcd;
8'hbe: tempout=8'h5a;
8'hbf: tempout=8'hf4;
8'hc0: tempout=8'h1f;
8'hc1: tempout=8'hdd;
8'hc2: tempout=8'ha8;
8'hc3: tempout=8'h33;
8'hc4: tempout=8'h88;
8'hc5: tempout=8'h07;
8'hc6: tempout=8'hc7;
8'hc7: tempout=8'h31;
8'hc8: tempout=8'hb1;
8'hc9: tempout=8'h12;
8'hca: tempout=8'h10;
8'hcb: tempout=8'h59;
8'hcc: tempout=8'h27;
8'hcd: tempout=8'h80;
8'hce: tempout=8'hec;
8'hcf: tempout=8'h5f;
8'hd0: tempout=8'h60;
8'hd1: tempout=8'h51;
8'hd2: tempout=8'h7f;
8'hd3: tempout=8'ha9;
8'hd4: tempout=8'h19;
8'hd5: tempout=8'hb5;
8'hd6: tempout=8'h4a;
8'hd7: tempout=8'h0d;
8'hd8: tempout=8'h2d;
8'hd9: tempout=8'he5;
8'hda: tempout=8'h7a;
8'hdb: tempout=8'h9f;
8'hdc: tempout=8'h93;
8'hdd: tempout=8'hc9;
8'hde: tempout=8'h9c;
8'hdf: tempout=8'hef;
8'he0: tempout=8'ha0;
8'he1: tempout=8'he0;
8'he2: tempout=8'h3b;
8'he3: tempout=8'h4d;
8'he4: tempout=8'hae;
8'he5: tempout=8'h2a;
8'he6: tempout=8'hf5;
8'he7: tempout=8'hb0;
8'he8: tempout=8'hc8;
8'he9: tempout=8'heb;
8'hea: tempout=8'hbb;
8'heb: tempout=8'h3c;
8'hec: tempout=8'h83;
8'hed: tempout=8'h53;
8'hee: tempout=8'h99;
8'hef: tempout=8'h61;
8'hf0: tempout=8'h17;
8'hf1: tempout=8'h2b;
8'hf2: tempout=8'h04;
8'hf3: tempout=8'h7e;
8'hf4: tempout=8'hba;
8'hf5: tempout=8'h77;
8'hf6: tempout=8'hd6;
8'hf7: tempout=8'h26;
8'hf8: tempout=8'he1;
8'hf9: tempout=8'h69;
8'hfa: tempout=8'h14;
8'hfb: tempout=8'h63;
8'hfc: tempout=8'h55;
8'hfd: tempout=8'h21;
8'hfe: tempout=8'h0c;
8'hff: tempout=8'h7d;
endcase





end



endmodule 